C:\Users\karl\Documents\NuTube\Nutubemk1.cir
* File created from design "C:\Users\karl\Documents\NuTube\Nutubemk1.sch" using DesignSpark 20.0.3

Tube1 N0024 N0024 N0043 N0050 ???? 
R1 N0024 3V3 150 
R2 N0023 3V3 150 
R3 3V3 GND 22K 
R4 N0043 N0030 10K 
IC1 N0015 3V3 
J1 N0002 GND GND FC681465P 
L1 12V N0002 10uH 
C3 12V GND 100nF 
C4 3V3 GND 100uF 
C2 N0002 GND 100uF 
C5 12V GND 100uF 
R7 N0015 GND 620 
R8 3V3 N0015 1K 
C6 N0015 GND 100nF 
C1 N0076 N0042 1uF 
R9 N0042 N0043 10K 
R5 3V3 GND 22k 
R6 N0046 N0044 10K 
C7 N0050 N0068 1uF 
R11 N0050 12V 330K 
R12 N0049 12V 330K 
C8 12V GND 100nF 
R13 N0060 N0084 100k 
C9 N0089 N0060 1uF 
R14 N0062 GND 100k 
C10 N0060 N0062 100nF 
R10 N0068 N0046 200k 
J2 N0072 GND GND 0449332 
J4 N0076 GND GND 0449332 
D1 N0002 GND SB5100 
C11 12V GND 100uF 
R15 N0084 GND 10K 
Q1 N0049 12V N0089 NMOS 
R16 N0089 GND 10K 
R17 N0049 N0089 DNI 
R18 3V3 N0100 150 
LED1 N0100 GND LED 5MM RED 
C12 3V3 GND 100nF 

.tran 0 1m 0 20u
.options Vntol=1u Abstol=1p Reltol=1m
.temp 27



.end
